// tw_im LUT, W=17 bits (2's complement)
case (addr)
  0: tw_im = 17'sh00000;
  1: tw_im = 17'sh1FFCE;
  2: tw_im = 17'sh1FF9C;
  3: tw_im = 17'sh1FF6A;
  4: tw_im = 17'sh1FF38;
  5: tw_im = 17'sh1FF07;
  6: tw_im = 17'sh1FED7;
  7: tw_im = 17'sh1FEA7;
  8: tw_im = 17'sh1FE78;
  9: tw_im = 17'sh1FE4A;
  10: tw_im = 17'sh1FE1D;
  11: tw_im = 17'sh1FDF2;
  12: tw_im = 17'sh1FDC7;
  13: tw_im = 17'sh1FD9E;
  14: tw_im = 17'sh1FD76;
  15: tw_im = 17'sh1FD50;
  16: tw_im = 17'sh1FD2C;
  17: tw_im = 17'sh1FD09;
  18: tw_im = 17'sh1FCE8;
  19: tw_im = 17'sh1FCCA;
  20: tw_im = 17'sh1FCAD;
  21: tw_im = 17'sh1FC92;
  22: tw_im = 17'sh1FC79;
  23: tw_im = 17'sh1FC62;
  24: tw_im = 17'sh1FC4E;
  25: tw_im = 17'sh1FC3C;
  26: tw_im = 17'sh1FC2C;
  27: tw_im = 17'sh1FC1F;
  28: tw_im = 17'sh1FC14;
  29: tw_im = 17'sh1FC0B;
  30: tw_im = 17'sh1FC05;
  31: tw_im = 17'sh1FC01;
  32: tw_im = 17'sh1FC00;
  33: tw_im = 17'sh1FC01;
  34: tw_im = 17'sh1FC05;
  35: tw_im = 17'sh1FC0B;
  36: tw_im = 17'sh1FC14;
  37: tw_im = 17'sh1FC1F;
  38: tw_im = 17'sh1FC2C;
  39: tw_im = 17'sh1FC3C;
  40: tw_im = 17'sh1FC4E;
  41: tw_im = 17'sh1FC62;
  42: tw_im = 17'sh1FC79;
  43: tw_im = 17'sh1FC92;
  44: tw_im = 17'sh1FCAD;
  45: tw_im = 17'sh1FCCA;
  46: tw_im = 17'sh1FCE8;
  47: tw_im = 17'sh1FD09;
  48: tw_im = 17'sh1FD2C;
  49: tw_im = 17'sh1FD50;
  50: tw_im = 17'sh1FD76;
  51: tw_im = 17'sh1FD9E;
  52: tw_im = 17'sh1FDC7;
  53: tw_im = 17'sh1FDF2;
  54: tw_im = 17'sh1FE1D;
  55: tw_im = 17'sh1FE4A;
  56: tw_im = 17'sh1FE78;
  57: tw_im = 17'sh1FEA7;
  58: tw_im = 17'sh1FED7;
  59: tw_im = 17'sh1FF07;
  60: tw_im = 17'sh1FF38;
  61: tw_im = 17'sh1FF6A;
  62: tw_im = 17'sh1FF9C;
  63: tw_im = 17'sh1FFCE;
  default: tw_im = '0;
endcase
