// tw_re LUT, W=17 bits (2's complement)
case (addr)
  0: tw_re = 17'sh00400;
  1: tw_re = 17'sh003FF;
  2: tw_re = 17'sh003FB;
  3: tw_re = 17'sh003F5;
  4: tw_re = 17'sh003EC;
  5: tw_re = 17'sh003E1;
  6: tw_re = 17'sh003D4;
  7: tw_re = 17'sh003C4;
  8: tw_re = 17'sh003B2;
  9: tw_re = 17'sh0039E;
  10: tw_re = 17'sh00387;
  11: tw_re = 17'sh0036E;
  12: tw_re = 17'sh00353;
  13: tw_re = 17'sh00336;
  14: tw_re = 17'sh00318;
  15: tw_re = 17'sh002F7;
  16: tw_re = 17'sh002D4;
  17: tw_re = 17'sh002B0;
  18: tw_re = 17'sh0028A;
  19: tw_re = 17'sh00262;
  20: tw_re = 17'sh00239;
  21: tw_re = 17'sh0020E;
  22: tw_re = 17'sh001E3;
  23: tw_re = 17'sh001B6;
  24: tw_re = 17'sh00188;
  25: tw_re = 17'sh00159;
  26: tw_re = 17'sh00129;
  27: tw_re = 17'sh000F9;
  28: tw_re = 17'sh000C8;
  29: tw_re = 17'sh00096;
  30: tw_re = 17'sh00064;
  31: tw_re = 17'sh00032;
  32: tw_re = 17'sh00000;
  33: tw_re = 17'sh1FFCE;
  34: tw_re = 17'sh1FF9C;
  35: tw_re = 17'sh1FF6A;
  36: tw_re = 17'sh1FF38;
  37: tw_re = 17'sh1FF07;
  38: tw_re = 17'sh1FED7;
  39: tw_re = 17'sh1FEA7;
  40: tw_re = 17'sh1FE78;
  41: tw_re = 17'sh1FE4A;
  42: tw_re = 17'sh1FE1D;
  43: tw_re = 17'sh1FDF2;
  44: tw_re = 17'sh1FDC7;
  45: tw_re = 17'sh1FD9E;
  46: tw_re = 17'sh1FD76;
  47: tw_re = 17'sh1FD50;
  48: tw_re = 17'sh1FD2C;
  49: tw_re = 17'sh1FD09;
  50: tw_re = 17'sh1FCE8;
  51: tw_re = 17'sh1FCCA;
  52: tw_re = 17'sh1FCAD;
  53: tw_re = 17'sh1FC92;
  54: tw_re = 17'sh1FC79;
  55: tw_re = 17'sh1FC62;
  56: tw_re = 17'sh1FC4E;
  57: tw_re = 17'sh1FC3C;
  58: tw_re = 17'sh1FC2C;
  59: tw_re = 17'sh1FC1F;
  60: tw_re = 17'sh1FC14;
  61: tw_re = 17'sh1FC0B;
  62: tw_re = 17'sh1FC05;
  63: tw_re = 17'sh1FC01;
  default: tw_re = '0;
endcase
